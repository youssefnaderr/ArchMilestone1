`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/10/2025 10:18:51 AM
// Design Name: 
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstMem (input [5:0] addr, output [31:0] data_out);

reg [31:0] mem[63:0];
assign data_out = mem[addr];
 
//R Type

//initial begin
//mem[0]= 32'b000000000101_00000_000_00010_0010011;  // ADDI x2, x0, 5
//mem[1]= 32'b000000000111_00000_000_00011_0010011; // ADDI x3, x0, 7
//mem[2]= 32'b0100000_00011_00010_000_00001_0110011;  // SUB x1, x2, x3
//mem[3]= 32'b0000000_00011_00010_001_00001_0110011;  // SLL x1, x2, x3
//mem[4]= 32'b0000000_00011_00010_010_00001_0110011;  // SLT x1, x2, x3
//mem[5]= 32'b0000000_00011_00010_011_00001_0110011;  // SLTU x1, x2, x3
//mem[6]= 32'b0000000_00011_00010_100_00001_0110011;  // XOR x1, x2, x3
//mem[7]= 32'b0000000_00011_00010_101_00001_0110011;  // SRL x1, x2, x3
//mem[8]= 32'b0100000_00011_00010_101_00001_0110011;  // SRA x1, x2, x3
//mem[9]= 32'b0000000_00011_00010_000_00001_0110011;  // ADD x1, x2, x3
//mem[10]= 32'b0000000_00011_00010_110_00001_0110011;  // OR x1, x2, x3
//mem[11]= 32'b0000000_00011_00010_111_00001_0110011;  // AND x1, x2, x3
//mem[12]= 32'b1111111_111111_11111_00001_1101111;  // JAL x1, -4
//end


//I Type

//initial begin
//mem[0] = 32'b000000000101_00000_000_00010_0010011;   // ADDI x2, x0, 5      
//mem[1] = 32'b0000000_00101_00010_001_00001_0010011;   // SLLI x1, x2, 5    
//mem[2] = 32'b000000001111_00010_010_00001_0010011;   // SLTI x1, x2, 15       
//mem[3] = 32'b0100000_00101_00010_101_00001_0010011;   // SRAI x1, x2, 5   
//mem[4] = 32'b0000000_00101_00010_101_00001_0010011;   // SRLI x1, x2, 5       
//mem[5] = 32'b000000000011_00010_011_00001_0010011;   // SLTIU x1, x2, 3      
//mem[6] = 32'b010000101010_00010_100_00001_0010011;   // XORI x1, x2, 42       
//mem[7] = 32'b000000010000_00010_110_00001_0010011;   // ORI x1, x2, 16        
//mem[8] = 32'b000000000111_00010_111_00001_0010011;   // ANDI x1, x2, 7       
//mem[9] = 32'b000000100000_00000_000_00000_1100111;   // JALR x0, 32(x0)    
//end


// BEQ
//initial begin
//mem[0] = 32'b000000000101_00000_000_00010_0010011 ;  // ADDI x2, x0, 5
//mem[1] = 32'b000000000101_00000_000_00011_0010011 ;  // ADDI x3, x0, 5
//mem[2] = 32'b0000000_00011_00010_000_00010_1100011 ; // BEQ x2, x3, +8
//mem[3] = 32'b0000000_00000_00000_000_00110_0110011 ; // ADD x6, x0, x0   (should be skipped)
//end

// BLT 

//initial begin
//mem[0] = 32'b000000000101_00000_000_00010_0010011 ;  // ADDI x2, x0, 5
//mem[1] = 32'b000000000110_00000_000_00011_0010011 ;  // ADDI x3, x0, 6
//mem[2] = 32'b0000000_00011_00010_100_00010_1100011 ; // BLT x2, x3, +8
//mem[3] = 32'b0000000_00000_00000_000_01000_0110011 ; // ADD x8, x0, x0   (should be skipped)
//end

// BGE

//initial
//mem[0] = 32'b000000000101_00000_000_00010_0010011 ;  // ADDI x2, x0, 5
//mem[1] = 32'b000000000100_00000_000_00011_0010011 ;  // ADDI x3, x0, 4
//mem[2] = 32'b0000000_00011_00010_101_00010_1100011 ; // BGE x2, x3, +8
//mem[3] = 32'b0000000_00000_00000_000_01001_0110011 ; // ADD x9, x0, x0   (should be skipped)
//end

// BLTU 

//initial
//mem[0] = 32'b000000000101_00000_000_00010_0010011 ;  // ADDI x2, x0, 5
//mem[1] = 32'b000000000110_00000_000_00011_0010011 ;  // ADDI x3, x0, 6
//mem[2] = 32'b0000000_00011_00010_110_00010_1100011 ; // BLTU x2, x3, +8
//mem[3] = 32'b0000000_00000_00000_000_01010_0110011 ; // ADD x10, x0, x0  (should be skipped)
//end

// BGEU 

//initial
//mem[0] = 32'b000000000101_00000_000_00010_0010011 ;  // ADDI x2, x0, 5
//mem[1] = 32'b000000000101_00000_000_00011_0010011 ;  // ADDI x3, x0, 5
//mem[2] = 32'b0000000_00011_00010_111_00010_1100011 ; // BGEU x2, x3, +8
//mem[3] = 32'b0000000_00000_00000_000_01011_0110011 ; // ADD x11, x0, x0  (should be skipped)
//end

// Load & PAUSE


//initial begin
//mem[0]= 32'b000000000000_00010_000_00001_0000011 ; // LB x1, 0(x2)
//mem[1]= 32'b000000000000_00010_001_00001_0000011;  // LH x1, 0(x2)
//mem[2]= 32'b000000000000_00010_010_00001_0000011;  // LW x1, 0(x2)
//mem[3]= 32'b000000000000_00010_100_00001_0000011;  // LBU x1, 0(x2)
//mem[4]= 32'b000000000000_00010_101_00001_0000011;  // LHU x1, 0(x2)  
//mem[5]= 32'b00000000000000000000000000001111;  // PAUSE
//end




//Store & LUI & AUIPC & ==EBREAK==


//initial begin
//mem[0]= 32'b000001111111_00000_000_00010_0010011 ;  // ADDI x2, x0, 2047
//mem[1]= 32'b000000001010_00000_000_00011_0010011;  // ADDI x3, x0, 10  
//mem[2] = 32'b0000000_00010_00000_010_00010_0100011 ; // SW x2, 2(x0)
//mem[3] = 32'b0000000_00010_00000_000_00010_0100011 ; // SB x2, 2(x0)
//mem[4] = 32'b0000000_00010_00000_001_00010_0100011 ; // SH x2, 2(x0)
//mem[5]= 32'b00010000000000000000_00001_0110111;  // LUI x1, 0x10000
//mem[6]= 32'b00010000000000000000_00001_0010111;  // AUIPC x1, 0x10000
//mem[7]= 32'b000000000001_00000_000_00000_1110011;  // EBREAK
//end


//Store & LUI & AUIPC & ==FENCE.TSO==

//initial begin
//mem[0]= 32'b000001111111_00000_000_00010_0010011 ;  // ADDI x2, x0, 2047
//mem[1]= 32'b000000001010_00000_000_00011_0010011;  // ADDI x3, x0, 10  
//mem[2] = 32'b0000000_00010_00000_010_00010_0100011 ; // SW x2, 2(x0)
//mem[3] = 32'b0000000_00010_00000_000_00010_0100011 ; // SB x2, 2(x0)
//mem[4] = 32'b0000000_00010_00000_001_00010_0100011 ; // SH x2, 2(x0)
//mem[5]= 32'b00010000000000000000_00001_0110111;  // LUI x1, 0x10000
//mem[6]= 32'b00010000000000000000_00001_0010111;  // AUIPC x1, 0x10000
//mem[7]= 32'b00001011000000000000000000001111;  // FENCE.TSO
//end


//Store & LUI & AUIPC & ==ECALL==


//initial begin
//mem[0]= 32'b000001111111_00000_000_00010_0010011 ;  // ADDI x2, x0, 2047
//mem[1]= 32'b000000001010_00000_000_00011_0010011;  // ADDI x3, x0, 10  
//mem[2] = 32'b0000000_00010_00000_010_00010_0100011 ; // SW x2, 2(x0)
//mem[3] = 32'b0000000_00010_00000_000_00010_0100011 ; // SB x2, 2(x0)
//mem[4] = 32'b0000000_00010_00000_001_00010_0100011 ; // SH x2, 2(x0)
//mem[5]= 32'b00010000000000000000_00001_0110111;  // LUI x1, 0x10000
//mem[6]= 32'b00010000000000000000_00001_0010111;  // AUIPC x1, 0x10000
//mem[7]= 32'b000000000000_00000_000_00000_1110011  // ECALL
//end



endmodule

